// Made by Aidan Ruck

MODULE maxJoltage;
ENDMODULE maxJoltage;
// This implementation (SystemVerilog instead of Verilog) does not need a module or package file, this is essentially here for show.